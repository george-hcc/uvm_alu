class environment extends uvm_environment;